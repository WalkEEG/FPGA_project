`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   09:09:14 07/27/2009
// Design Name:   epinout
// Module Name:   E:/ZYQ/work/ISE/usb/UART/adfifo/fifotestf.v
// Project Name:  adfifotest
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: epinout
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module processtest;

	 reg clk = 1'b0;
	 reg clk1_2 =1'b0;
    reg en = 1'b0;
	 reg reset =1'b0;
    reg ad_clk = 1'b0;
    reg ad_data = 1'b0;
	 reg ad_ready = 1'b0;
	 
	 reg syn_head_tb1 = 1'b0;
	 reg syn_head_tb2 = 1'b0;
    wire [7:0]ramdata;
	 
    parameter PERIOD = 100;
    parameter real DUTY_CYCLE = 0.5;
    parameter OFFSET = 50;

    initial    // Clock process for clk
    begin
        #OFFSET;
        forever
        begin
            clk = 1'b0;
				#(PERIOD-(PERIOD*DUTY_CYCLE)) clk = 1'b1;
            #(PERIOD*DUTY_CYCLE);
		  end
    end
	 
initial    // Clock process for clk
    begin
        #OFFSET;
        forever
        begin
            clk1_2 = 1'b0;
				#25 clk1_2 = 1'b1;
            #25;
		  end
    end

	///
    processmain UUT (
        .clk(clk),
		  .clk1_2(clk1_2),
        .en(en),
		  .reset(reset),
		  
		  .ad_clk(ad_clk),       
        .ad_data(ad_data),
		  .ad_ready(ad_ready),
		  
		  .syn_head_tb1(syn_head_tb1),
		  .syn_head_tb2(syn_head_tb2),
		  .ramdata(ramdata)		  
		  );

    initial begin
        // -------------  Current Time:  185ns
      
        en = 1'b1;
		  reset=1'b1;
        // -------------------------------------
        // -------------  Current Time:  1185ns
 forever
        begin
		  
        #100;
		  ad_ready=1;
		  #100;
		  ad_ready=0;
		  
		  #100;
        ad_clk = 1'b1;
		  ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  6185ns
        #100;
        ad_clk = 1'b0;
		  ad_data= 1'b0;
//ad_count==1		  
        // -------------------------------------
        // -------------  Current Time:  11185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  16185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==2		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==3
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==4		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==5
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==6		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==7
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;	
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1; 
//ad_count==8		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==9
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;

//ad_count==10
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==11		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==12
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;		  

//ad_count==13
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==14		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==15
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==16		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==17
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
		  
//ad_count==18
		  #100;
		  ad_clk = 1'b1;
		  ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  6185ns
        #100;
        ad_clk = 1'b0;
		  ad_data= 1'b1;
//ad_count==19		  
        // -------------------------------------
        // -------------  Current Time:  11185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  16185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==20		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==21
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==22		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==23
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==0		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
		  
//ad_count==1
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;	
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0; 
//ad_count==2		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==3
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;

//ad_count==4
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==5		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==6
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;		  

//ad_count==7
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==8		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==9
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==10		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==11
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
	
//ad_count==12
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;		  

//ad_count==13
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==14		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==15
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==16		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==17
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
		  
//ad_count==18
		  #100;
		  ad_clk = 1'b1;
		  ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  6185ns
        #100;
        ad_clk = 1'b0;
		  ad_data= 1'b0;
//ad_count==19		  
        // -------------------------------------
        // -------------  Current Time:  11185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  16185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==20		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==21
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==22		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==23
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;	
		  
	//#1000;
//ad_count==0
		        #100;
        ad_clk = 1'b1;
		  ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  6185ns
        #100;
        ad_clk = 1'b0;
		  ad_data= 1'b1;
//ad_count==1		  
        // -------------------------------------
        // -------------  Current Time:  11185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  16185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==2		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==3
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==4		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==5
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==6		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==7
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;	
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1; 
//ad_count==8		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==9
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;

//ad_count==10
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==11		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==12
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;		  

//ad_count==13
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==14		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==15
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==16		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==17
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
		  
//ad_count==18
		  #100;
		  ad_clk = 1'b1;
		  ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  6185ns
        #100;
        ad_clk = 1'b0;
		  ad_data= 1'b1;
//ad_count==19		  
        // -------------------------------------
        // -------------  Current Time:  11185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  16185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==20		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==21
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==22		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==23
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==0		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
		  
//ad_count==1
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;	
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1; 
//ad_count==2		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==3
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;

//ad_count==4
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==5		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==6
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;		  

//ad_count==7
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==8		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==9
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==10		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==11
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
	
//ad_count==12
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;		  

//ad_count==13
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==14		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==15
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==16		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==17
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
		  
//ad_count==18
		  #100;
		  ad_clk = 1'b1;
		  ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  6185ns
        #100;
        ad_clk = 1'b0;
		  ad_data= 1'b1;
//ad_count==19		  
        // -------------------------------------
        // -------------  Current Time:  11185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  16185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==20		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==21
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==22		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==23
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;	
        // -------------  Current Time:  1185ns
        #100;
        ad_clk = 1'b1;
		  ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  6185ns
        #100;
        ad_clk = 1'b0;
		  ad_data= 1'b0;
//ad_count==1		  
        // -------------------------------------
        // -------------  Current Time:  11185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  16185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==2		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==3
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==4		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==5
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==6		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==7
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;	
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1; 
//ad_count==8		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==9
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;

//ad_count==10
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==11		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==12
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;		  

//ad_count==13
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==14		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==15
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==16		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==17
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
		  
//ad_count==18
		  #100;
		  ad_clk = 1'b1;
		  ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  6185ns
        #100;
        ad_clk = 1'b0;
		  ad_data= 1'b1;
//ad_count==19		  
        // -------------------------------------
        // -------------  Current Time:  11185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  16185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==20		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==21
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==22		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==23
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b1;
//ad_count==0		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
		  
//ad_count==1
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;	
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0; 
//ad_count==2		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==3
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;

//ad_count==4
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==5		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==6
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;		  

//ad_count==7
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==8		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==9
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==10		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==11
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
	
//ad_count==12
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;		  

//ad_count==13
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==14		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==15
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==16		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==17
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
		  
//ad_count==18
		  #100;
		  ad_clk = 1'b1;
		  ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  6185ns
        #100;
        ad_clk = 1'b0;
		  ad_data= 1'b0;
//ad_count==19		  
        // -------------------------------------
        // -------------  Current Time:  11185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  16185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==20		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==21
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data =1'b0;
//ad_count==22		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==23
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;	
		  
	//#1000;
//ad_count==0
		        #100;
        ad_clk = 1'b1;
		  ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  6185ns
        #100;
        ad_clk = 1'b0;
		  ad_data= 1'b1;
//ad_count==1		  
        // -------------------------------------
        // -------------  Current Time:  11185ns
        #100;
        ad_clk = 1'b1;
        ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  16185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==2		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==3
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==4		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==5
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==6		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==7
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;	
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1; 
//ad_count==8		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==9
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;

//ad_count==10
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==11		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==12
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;		  

//ad_count==13
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==14		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==15
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==16		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==17
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
		  
//ad_count==18
		  #100;
		  ad_clk = 1'b1;
		  ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  6185ns
        #100;
        ad_clk = 1'b0;
		  ad_data= 1'b1;
//ad_count==19		  
        // -------------------------------------
        // -------------  Current Time:  11185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  16185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==20		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==21
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==22		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==23
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==0		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
		  
//ad_count==1
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;	
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1; 
//ad_count==2		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==3
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;

//ad_count==4
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==5		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==6
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;		  

//ad_count==7
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==8		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==9
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==10		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==11
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
	
//ad_count==12
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;		  

//ad_count==13
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==14		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==15
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==16		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==17
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
		  
//ad_count==18
		  #100;
		  ad_clk = 1'b1;
		  ad_data =1'b1;
        // -------------------------------------
        // -------------  Current Time:  6185ns
        #100;
        ad_clk = 1'b0;
		  ad_data= 1'b1;
//ad_count==19		  
        // -------------------------------------
        // -------------  Current Time:  11185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  16185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==20		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==21
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;
//ad_count==22		 
		  // -------------------------------------
        // -------------  Current Time:  21185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b0;
        // -------------------------------------
        // -------------  Current Time:  26185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b0;
//ad_count==23
        // -------------------------------------
        // -------------  Current Time:  31185ns
        #100;
        ad_clk = 1'b1;
        ad_data = 1'b1;
        // -------------------------------------
        // -------------  Current Time:  36185ns
        #100;
        ad_clk = 1'b0;
        ad_data = 1'b1;	
		  
		  #1000;
		  end
	 end

      
endmodule

